*******************************************************************************
* CDL netlist
*
* Library : New_lib
* Top Cell Name: aoi
* View Name: layout
* Netlist created: 4.Jul.2017
*******************************************************************************

*.SCALE METER
*.GLOBAL 

*******************************************************************************
* Library Name: New_lib
* Cell Name:    aoi
* View Name:    layout
*******************************************************************************

.SUBCKT aoi
*.PININFO

.ENDS
