*******************************************************************************
* CDL netlist
*
* Library : NangateOpenCellLibrary
* Top Cell Name: Nand
* View Name: layout
* Netlist created: 7.Jul.2017
*******************************************************************************

*.SCALE METER
*.GLOBAL addEnd 0 

*******************************************************************************
* Library Name: NangateOpenCellLibrary
* Cell Name:    Nand
* View Name:    layout
*******************************************************************************

.SUBCKT Nand

.ENDS
