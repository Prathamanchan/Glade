   /   0   
Inverter2    1   
extracted    2   3   I  �   J>.�&֕   K          x   �  ;             �      text       drawing          �        M1                 ?�         F       A         �  �      M0                 ?�         F       A   A          POLY       drawing          Y  	�    	�    �  �  �  �  	�  �  	�  �  h  �  h  �  �    �    h  Y  h      n2    A   A    	      NIMP       drawing         d      �      n4    A        	�  �  ~  �      n5    A   A           PWELL       drawing         �  q  6  
K      n0    A   A    
      CONT       drawing         �  �  �  u      n1    A        �  �  �  �      n1    A        �  �  �  �      n1    A        �  �  �  �      n1    A        �    �  �      n1    A        �  &  �        n0    A        �  F  �  "      n0    A        �  �  �  u      n1    A        �  �  �  �      n1    A        �  �  �  �      n1    A        �    �  �      n1    A        �  
  �  
�      n2    A        �  �  �  �      n1    A        �  F  �  "      n0    A        �  &  �        n0    A        �  
  ~  
�      n2    A        �  �  �  u      n3    A        �  �  �  �      n3    A        �  �  �  �      n3    A        �    �  �      n3    A        �  �  �  �      n3    A        �  F  �  "      n3    A        �  &  �        n3    A   A          DIFF       drawing         �  *  ~  �      n3    A        	�  *    �      n1    A        d  �    z      n0    A        d      �      n1    A        	�  �    �      n0    A        �  �  ~  �      n3    A   A   �      	instance       drawing            *          D?�                  M1       PCH_SVT_1P8V_EX       layout        *  �  �                !       "             w    	      G   
>�*sq�T      l    	      G   
>�/��߸      as    	      G   
=��{��6      ps    	      G   
>��u�Nj      ad    	      G   
=��J��      pd    	      G   
>���k�   4      &   B       n1    (    &   D       n3    (    &   S       n1    (    &   G       n2    (    A           �          D?�                  M0       NCH_SVT_1P8V_EX       layout        �  �  �                !       "             w    	      G   
>������      l    	      G   
>�/��߸      as    	      G   
=sY����y      ps    	      G   
>��򚼯H      ad    	      G   
=q=�ec      pd    	      G   
>�ԍ5�"$   4      &   B       n0    (    &   D       n3    (    &   S       n0    (    &   G       n2    (    A   A          MET1       drawing           x  ]    ]    b  _  b  _            b  �  b  �  9  �  9  �  b  �  b  �  �  �  �  �    �    �  �   x  �      n1    A            �  d   �  d    �    �  �  �  �  �          p  i  p  i    �    �  !    !              n0    A        	t  	�  A  h      n2    A        �  �  �  �      n3    A   A          PIMP       drawing         d  �    z      n6    A        	�  *  ~  �      n7    A   A          NWELL       drawing         �  J  ;  �      n1    A   A   4      n6    )    5          n1    )    5          n3    )    5          n4    )    5          n0    )    5          n2    )    5          n7    )    5          n5    )    5       A